library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TRIANGLE_WAVE_GEN is
	port(
		CLK, INV: in std_logic;
		wave : out std_logic_vector(7 downto 0)
	);
end entity;

architecture func of TRIANGLE_WAVE_GEN is
	
	begin
--	--======================================================================================================================--
--	process(CLK) begin
--
--	end process;
	
end architecture;