library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity COUNTER_3_BITS is
	port(
		CLK : in std_logic;
		C : out std_logic_vector(2 downto 0)
	);
end entity;

architecture count of COUNTER_3_BITS is
begin
	--
end architecture;