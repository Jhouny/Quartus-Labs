library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity COMPARATOR_8_BITS is
	port(
		A, REF : in std_logic_vector(7 downto 0);
		Q : out std_logic
	);
end entity;

architecture func of COMPARATOR_8_BITS is
	begin
end architecture;