library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SQUARE_WAVE_GEN_50 is
	port(
		COUNT: in std_logic_vector(7 downto 0);
		wave : out std_logic_vector(7 downto 0)
	);
end entity;

architecture func of SQUARE_WAVE_GEN_50 is
	
	begin
--	--======================================================================================================================--
--	process(CLK) begin
--
--	end process;
	
end architecture;